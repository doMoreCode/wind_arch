module Not(input in, output out);
  // your code here
  Nand g1(in, in, out);

endmodule



