module FullAdder(input a,b,c, output sum, carry);
  // your code here

endmodule
